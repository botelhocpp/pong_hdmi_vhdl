LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

PACKAGE HdmiPkg IS 
    SUBTYPE t_Byte IS STD_LOGIC_VECTOR(7 DOWNTO 0);
    SUBTYPE t_RGB IS STD_LOGIC_VECTOR(23 DOWNTO 0);
    
    CONSTANT c_FRAME_WIDTH   : INTEGER := 640;
    CONSTANT c_H_FRONT_PORCH : INTEGER := 16;
    CONSTANT c_H_BACK_PORCH  : INTEGER := 48;
    CONSTANT c_H_PULSE_WIDTH : INTEGER := 96;
    CONSTANT c_H_BLANK       : INTEGER := c_H_FRONT_PORCH + c_H_BACK_PORCH + c_H_PULSE_WIDTH;
    
    CONSTANT c_FRAME_HEIGHT    : INTEGER := 480;
    CONSTANT c_V_FRONT_PORCH   : INTEGER := 10;
    CONSTANT c_V_BACK_PORCH    : INTEGER := 33;
    CONSTANT c_V_PULSE_WIDTH   : INTEGER := 2;
    CONSTANT c_V_BLANK         : INTEGER := c_V_FRONT_PORCH + c_V_BACK_PORCH + c_V_PULSE_WIDTH;
    
    CONSTANT c_H_MAX : INTEGER := c_FRAME_WIDTH + c_H_BLANK;
    CONSTANT c_V_MAX : INTEGER := c_FRAME_HEIGHT + c_V_BLANK;
	
	CONSTANT c_DISPLAY_RESOLUTION : INTEGER := c_FRAME_WIDTH * c_FRAME_HEIGHT;
	CONSTANT c_MAX_RESOLUTION : INTEGER := c_H_MAX * c_V_MAX;  

END HdmiPkg;
