LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
 
LIBRARY WORK;
USE WORK.HdmiPkg.ALL;

PACKAGE PongPkg IS
  CONSTANT c_GAME_SCALE : INTEGER := 20;
  
  CONSTANT c_REFRESH_RATE : INTEGER := c_PIXEL_CLK_FREQ/c_GAME_SCALE;
  CONSTANT c_GAME_WIDTH : INTEGER := c_FRAME_WIDTH/c_GAME_SCALE;
  CONSTANT c_GAME_HEIGHT : INTEGER := c_FRAME_HEIGHT/c_GAME_SCALE;
 
  CONSTANT c_SCORE_LIMIT : INTEGER := 9;
  CONSTANT c_SCORE_WIDTH : INTEGER := 3;
  CONSTANT c_SCORE_HEIGHT : INTEGER := 5;
  CONSTANT c_SCORE_Y_POS : INTEGER := 1;
   
  CONSTANT c_PADDLE_HEIGHT : INTEGER := 6;
  
  CONSTANT c_PADDLE_SPEED : INTEGER := c_REFRESH_RATE; 
  CONSTANT c_BALL_SPEED : INTEGER  := c_REFRESH_RATE;
   
  CONSTANT c_P1_PADDLE_COL : INTEGER := 0;
  CONSTANT c_P2_PADDLE_COL : INTEGER := c_GAME_WIDTH - 1;
  CONSTANT c_P1_SCORE_COL : INTEGER := c_GAME_WIDTH/2 - 2*c_SCORE_WIDTH - c_SCORE_WIDTH;
  CONSTANT c_P2_SCORE_COL : INTEGER := c_GAME_WIDTH/2 + 2*c_SCORE_WIDTH;
  
END PACKAGE PongPkg; 