LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
 
LIBRARY WORK;
USE WORK.HdmiPkg.ALL;

PACKAGE PongPkg IS
  CONSTANT c_GAME_WIDTH : INTEGER := c_FRAME_WIDTH/16;
  CONSTANT c_GAME_HEIGHT : INTEGER := c_FRAME_HEIGHT/16;
 
  CONSTANT c_SCORE_LIMIT : INTEGER := 9;
  CONSTANT c_SCORE_WIDTH : INTEGER := 3;
  CONSTANT c_SCORE_HEIGHT : INTEGER := 5;
  CONSTANT c_SCORE_Y_POS : INTEGER := 2;
   
  CONSTANT c_PADDLE_HEIGHT : INTEGER := 6;
 
  CONSTANT c_PADDLE_SPEED : INTEGER := 1250000; 
  CONSTANT c_BALL_SPEED : INTEGER  := 1250000;
   
  CONSTANT c_P1_PADDLE_COL : INTEGER := 0;
  CONSTANT c_P2_PADDLE_COL : INTEGER := c_GAME_WIDTH - 1;
  
END PACKAGE PongPkg; 